-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 12.1 Build 177 11/07/2012 SJ Full Version"
-- CREATED		"Fri Sep 13 15:05:34 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY prime2 IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC;
		E :  IN  STD_LOGIC;
		F :  IN  STD_LOGIC;
		O :  OUT  STD_LOGIC
	);
END prime2;

ARCHITECTURE bdf_type OF prime2 IS 

SIGNAL	o_ALTERA_SYNTHESIZED17 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED19 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED23 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED29 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED31 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED37 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED41 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED43 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED47 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED53 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED59 :  STD_LOGIC;
SIGNAL	o_ALTERA_SYNTHESIZED61 :  STD_LOGIC;
SIGNAL	prum :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;


BEGIN 



o_ALTERA_SYNTHESIZED17 <= SYNTHESIZED_WIRE_0 AND A AND SYNTHESIZED_WIRE_1 AND SYNTHESIZED_WIRE_2 AND E AND SYNTHESIZED_WIRE_3;


o_ALTERA_SYNTHESIZED19 <= SYNTHESIZED_WIRE_4 AND A AND B AND SYNTHESIZED_WIRE_5 AND E AND SYNTHESIZED_WIRE_6;


o_ALTERA_SYNTHESIZED23 <= C AND A AND B AND SYNTHESIZED_WIRE_7 AND E AND SYNTHESIZED_WIRE_8;


o_ALTERA_SYNTHESIZED29 <= C AND A AND SYNTHESIZED_WIRE_9 AND D AND E AND SYNTHESIZED_WIRE_10;


o_ALTERA_SYNTHESIZED31 <= C AND A AND B AND D AND E AND SYNTHESIZED_WIRE_11;


o_ALTERA_SYNTHESIZED37 <= C AND A AND SYNTHESIZED_WIRE_12 AND SYNTHESIZED_WIRE_13 AND SYNTHESIZED_WIRE_14 AND F;


o_ALTERA_SYNTHESIZED41 <= SYNTHESIZED_WIRE_15 AND A AND SYNTHESIZED_WIRE_16 AND D AND SYNTHESIZED_WIRE_17 AND F;


o_ALTERA_SYNTHESIZED43 <= SYNTHESIZED_WIRE_18 AND A AND B AND D AND SYNTHESIZED_WIRE_19 AND F;


o_ALTERA_SYNTHESIZED47 <= C AND A AND B AND D AND SYNTHESIZED_WIRE_20 AND F;


o_ALTERA_SYNTHESIZED53 <= C AND A AND SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_22 AND E AND F;


o_ALTERA_SYNTHESIZED59 <= SYNTHESIZED_WIRE_23 AND A AND B AND D AND E AND F;


o_ALTERA_SYNTHESIZED61 <= C AND A AND SYNTHESIZED_WIRE_24 AND D AND E AND F;


prum <= o_ALTERA_SYNTHESIZED23 OR o_ALTERA_SYNTHESIZED19 OR o_ALTERA_SYNTHESIZED17 OR o_ALTERA_SYNTHESIZED31 OR o_ALTERA_SYNTHESIZED47 OR o_ALTERA_SYNTHESIZED29 OR o_ALTERA_SYNTHESIZED41 OR o_ALTERA_SYNTHESIZED37 OR o_ALTERA_SYNTHESIZED43 OR o_ALTERA_SYNTHESIZED59 OR o_ALTERA_SYNTHESIZED53 OR o_ALTERA_SYNTHESIZED61;


SYNTHESIZED_WIRE_25 <= A AND B AND C AND D;


SYNTHESIZED_WIRE_33 <= NOT(SYNTHESIZED_WIRE_25);



SYNTHESIZED_WIRE_32 <= NOT(F);



SYNTHESIZED_WIRE_3 <= NOT(F);



SYNTHESIZED_WIRE_36 <= A AND SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_1 <= NOT(B);



SYNTHESIZED_WIRE_0 <= NOT(C);



SYNTHESIZED_WIRE_2 <= NOT(D);



SYNTHESIZED_WIRE_6 <= NOT(F);



SYNTHESIZED_WIRE_8 <= NOT(F);



SYNTHESIZED_WIRE_4 <= NOT(C);



SYNTHESIZED_WIRE_35 <= SYNTHESIZED_WIRE_27 AND B AND SYNTHESIZED_WIRE_28 AND SYNTHESIZED_WIRE_29;


SYNTHESIZED_WIRE_5 <= NOT(D);



SYNTHESIZED_WIRE_10 <= NOT(F);



SYNTHESIZED_WIRE_9 <= NOT(B);



SYNTHESIZED_WIRE_7 <= NOT(D);



SYNTHESIZED_WIRE_11 <= NOT(F);



SYNTHESIZED_WIRE_12 <= NOT(B);



SYNTHESIZED_WIRE_16 <= NOT(B);



SYNTHESIZED_WIRE_13 <= NOT(D);



SYNTHESIZED_WIRE_14 <= NOT(E);



SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_31 AND SYNTHESIZED_WIRE_32 AND SYNTHESIZED_WIRE_33;


SYNTHESIZED_WIRE_15 <= NOT(C);



SYNTHESIZED_WIRE_21 <= NOT(B);



SYNTHESIZED_WIRE_17 <= NOT(E);



SYNTHESIZED_WIRE_18 <= NOT(C);



SYNTHESIZED_WIRE_24 <= NOT(B);



SYNTHESIZED_WIRE_19 <= NOT(E);



SYNTHESIZED_WIRE_22 <= NOT(D);



SYNTHESIZED_WIRE_20 <= NOT(E);



SYNTHESIZED_WIRE_23 <= NOT(C);



SYNTHESIZED_WIRE_31 <= NOT(E);



O <= prum OR SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_26 <= C OR B;


SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_35 OR SYNTHESIZED_WIRE_36;


SYNTHESIZED_WIRE_27 <= NOT(A);



SYNTHESIZED_WIRE_28 <= NOT(C);



SYNTHESIZED_WIRE_29 <= NOT(D);



END bdf_type;