-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 12.1 Build 177 11/07/2012 SJ Full Version"
-- CREATED		"Tue Sep 10 12:25:49 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY traffic IS 
	PORT
	(
		enable :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		NSred :  OUT  STD_LOGIC;
		EWred :  OUT  STD_LOGIC;
		NSyellow :  OUT  STD_LOGIC;
		EWyellow :  OUT  STD_LOGIC;
		NSgreen :  OUT  STD_LOGIC;
		EWgreen :  OUT  STD_LOGIC;
		q :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END traffic;

ARCHITECTURE bdf_type OF traffic IS 

COMPONENT counter
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 enable : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	q_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_4 <= '1';



SYNTHESIZED_WIRE_2 <= q_ALTERA_SYNTHESIZED(2) XOR q_ALTERA_SYNTHESIZED(1);


EWred <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3;


b2v_inst : counter
PORT MAP(clk => clk,
		 reset => reset,
		 enable => SYNTHESIZED_WIRE_4,
		 q => q_ALTERA_SYNTHESIZED);


SYNTHESIZED_WIRE_11 <= SYNTHESIZED_WIRE_5 AND SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_7;


SYNTHESIZED_WIRE_1 <= NOT(q_ALTERA_SYNTHESIZED(3));



SYNTHESIZED_WIRE_0 <= q_ALTERA_SYNTHESIZED(3) AND SYNTHESIZED_WIRE_8 AND SYNTHESIZED_WIRE_9 AND SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_21 <= NOT(SYNTHESIZED_WIRE_11);



SYNTHESIZED_WIRE_8 <= NOT(q_ALTERA_SYNTHESIZED(2));



SYNTHESIZED_WIRE_9 <= NOT(q_ALTERA_SYNTHESIZED(1));



SYNTHESIZED_WIRE_10 <= NOT(q_ALTERA_SYNTHESIZED(0));



SYNTHESIZED_WIRE_6 <= NOT(q_ALTERA_SYNTHESIZED(1));



SYNTHESIZED_WIRE_7 <= NOT(q_ALTERA_SYNTHESIZED(0));




SYNTHESIZED_WIRE_3 <= q_ALTERA_SYNTHESIZED(0) AND SYNTHESIZED_WIRE_12 AND SYNTHESIZED_WIRE_13;


SYNTHESIZED_WIRE_12 <= NOT(q_ALTERA_SYNTHESIZED(1));



SYNTHESIZED_WIRE_13 <= NOT(q_ALTERA_SYNTHESIZED(2));



NSgreen <= SYNTHESIZED_WIRE_14 AND SYNTHESIZED_WIRE_15;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_16 AND SYNTHESIZED_WIRE_17 AND SYNTHESIZED_WIRE_18 AND SYNTHESIZED_WIRE_19;


SYNTHESIZED_WIRE_16 <= NOT(q_ALTERA_SYNTHESIZED(3));



SYNTHESIZED_WIRE_17 <= NOT(q_ALTERA_SYNTHESIZED(2));



SYNTHESIZED_WIRE_18 <= NOT(q_ALTERA_SYNTHESIZED(1));



SYNTHESIZED_WIRE_19 <= NOT(q_ALTERA_SYNTHESIZED(0));



SYNTHESIZED_WIRE_14 <= NOT(q_ALTERA_SYNTHESIZED(3));



EWgreen <= q_ALTERA_SYNTHESIZED(3) AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21;


NSred <= SYNTHESIZED_WIRE_22 OR q_ALTERA_SYNTHESIZED(3);


NSyellow <= SYNTHESIZED_WIRE_23 AND q_ALTERA_SYNTHESIZED(2) AND q_ALTERA_SYNTHESIZED(1);


SYNTHESIZED_WIRE_5 <= NOT(q_ALTERA_SYNTHESIZED(2));



SYNTHESIZED_WIRE_23 <= NOT(q_ALTERA_SYNTHESIZED(3));



EWyellow <= q_ALTERA_SYNTHESIZED(3) AND q_ALTERA_SYNTHESIZED(2) AND q_ALTERA_SYNTHESIZED(1);


SYNTHESIZED_WIRE_20 <= NOT(q_ALTERA_SYNTHESIZED(1) AND q_ALTERA_SYNTHESIZED(2));

q <= q_ALTERA_SYNTHESIZED;

END bdf_type;